`include "uvm_pkg.sv"
import uvm_pkg::*;
`include "usbf_defines.v"
`include "usbf_crc16.v"
`include "usbf_crc5.v"
`include "usbf_ep_rf_dummy.v"
`include "usbf_ep_rf.v"
`include "usbf_idma.v"
`include "usbf_mem_arb.v"
`include "usbf_pa.v"
`include "usbf_pd.v"
`include "usbf_pe.v"
`include "usbf_pl.v"
`include "usbf_rf.v"
`include "usbf_utmi_if.v"
`include "usbf_utmi_ls.v"
`include "usbf_wb.v"
`include "usbf_top.v"
`include "utmi_intf.sv"
`include "wb_intf.sv"
`include "wb_tx.sv"
`include "reg2wb_adapter.sv"
`include "usb_reg_model.sv"
`include "usb_config.sv"
`include "wb_sequence_lib.sv"
`include "usb_frame.sv"
`include "utmi_sequence_lib.sv"
`include "utmi_driver.sv"
`include "utmi_sqr.sv"
`include "utmi_mon.sv"
`include "utmi_cov.sv"
`include "utmi_agent.sv"
`include "wb_cov.sv"
`include "wb_sqr.sv"
`include "wb_driver.sv"
`include "wb_mon.sv"
`include "wb_agent.sv"
`include "usb_sbd.sv"
`include "usb_top_sqr.sv"
`include "usb_seq_lib.sv"
`include "usb_env.sv"
`include "top.sv"
